
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity task3 is
    Port (
        sw  : in  std_logic_vector(15 downto 0);  -- ���������� ������� 8 ���
        led : out std_logic_vector(15 downto 0)
    );
end task3;
--������� 5 K = 31B6(16) = 11 0001 1011 0110(2) = 14 ��� I = D5 J = 7A F = 31B6 A = and B = + C = >>3 D = nor G = ���� (7 ���) L = 6420
architecture Behavioral of task3 is
    constant I : std_logic_vector(7 downto 0) := x"D5"; -- 11010101
    constant J : std_logic_vector(7 downto 0) := x"7A"; -- 01111010
begin

    -- ������ ��������: led_o[7:0] = sw_i[7:0] XOR I
    led(7 downto 0) <= sw(7 downto 0) xor I     ;

    -- ��������� ���� J, ����� ��� 16 LED ���?�� ����������:
    led(15 downto 8) <= J;  -- ��������, ��������� J �� ������� 8 �����������

end Behavioral;
